//Define all characters with the 4bit value
//Author Tselepi Eleni 03272

`define zero 4'b0000
`define one 4'b0001
`define two 4'b0010
`define three 4'b0011
`define four 4'b0100
`define five 4'b0101
`define six 4'b0110
`define seven 4'b0111
`define eight 4'b1000
`define nine 4'b1001
`define a 4'b1010
`define b 4'b1011
`define c 4'b1100
`define d 4'b1101
`define e 4'b1110
`define F 4'b1111