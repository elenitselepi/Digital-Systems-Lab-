//Define all time distances in cycles for the hsync

`define A 'd3200
`define B 'd384
`define C 'd192
`define D 'd2560
`define E 'd64