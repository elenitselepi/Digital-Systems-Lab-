//Define all time distances in cycles for vsync

`define O 'd1_667_200
`define P 'd6400
`define Q 'd92_800
`define R 'd1_536_000
`define S 'd32_000